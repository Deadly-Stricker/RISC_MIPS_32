module IF_stage(
    input clk,
    input stall,
    input [31:0]Next_pc,
    input jump_cs,
    output reg [31:0]instruction
);
    wire connector_from_pc_to_IR; 
    // reg Instruction_storage;
    programCounter PC_Module (.clk(clk),.stall(stall),.Next_pc(Next_pc),.jump_cs(jump_cs),.pc_curr(connector_from_pc_to_IR));
    instructionRegister IR_Module (.clk(clk),.pc(connector_from_pc_to_IR),.instruction(instruction));

endmodule